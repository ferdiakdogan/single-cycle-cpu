module instruction_memory #(parameter ADDR_WIDTH = 32, DATA_WIDTH = 32) (
	in, out
);

	input [ADDR_WIDTH-1:0] in;
	output [DATA_WIDTH-1:0] out;

	reg [DATA_WIDTH-1:0] memory [127:0];
	
	initial begin
		memory [0] = 32'b11100010100000010001000000000010; //r1 = 2
		memory [4] = 32'b11100010100000100010000000000011; //r2 = 3
		memory [8] = 32'b11100010100000110011000000000100; //r3 = 4
		memory [12] = 32'b11100010100001000100000000000101; //r4 = 5
		memory [16] = 32'b11100010100001010101000000000110; //r5 = 6
		memory [20] = 32'b11100010100001100110000000000111; //r6 = 7
		memory [24] = 32'b11100010100001110111000000001000; //r7 = 8
		memory [28] = 32'b11100010100010001000000000001001; //r8 = 9
		memory [32] = 32'b11100000100000010000000000000010; //r0 = r1+r2
		memory [36] = 32'b11100000010001110000000000000100; //r0 = r7 - r4
		memory [40] = 32'b11100000000000000000000000000001; // r0 = r0 & r1
		memory [44] = 32'b11100001100000000000000000000010; // r0 = r0 | r1
		memory [48] = 32'b11100001101000000000000010100000; // lsr r0, r0, #1
		memory [52] = 32'b11100001101000000000000100000000; // lsl r0, r0, #2
		memory [56] = 32'b11100001010100110000000000000000; // cmp r0, r3
		memory [60] = 32'b11100101101000010110000000000110; // str r6,[r1,#6]
		memory [64] = 32'b11100101100100010000000000000110; // ldr r0,[r1,#6]
	end
	
	
	assign out = memory[in];
	
endmodule